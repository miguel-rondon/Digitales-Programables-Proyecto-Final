LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY LIB_TEC_MATRICIAL_4x4_INTESC_RevA IS
	--El generic es útil cuando LIB_TEC_MATRICIAL_4x4_INTESC_RevA es parte de un TOP. Si no es parte de un TOP
	--entonces se deben poner la frecuencia del FPGA como valores contantes en el generic
	GENERIC (
		FREQ_CLK : INTEGER := 50_000_000 --FRECUENCIA DE LA TARJETA
	);
	PORT (
		CLK : IN STD_LOGIC; --RELOJ FPGA
		COLUMNAS : IN STD_LOGIC_VECTOR(3 DOWNTO 0); --PUERTO CONECTADO A LAS COLUMNAS DEL TECLADO
		FILAS : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); --PUERTO CONECTADO A LA FILAS DEL TECLADO
		BOTON_PRES : OUT STD_LOGIC_VECTOR(3 DOWNTO 0); --PUERTO QUE INDICA LA TECLA QUE SE PRESIONÓ
		IND : OUT STD_LOGIC --BANDERA QUE INDICA CUANDO SE PRESIONÓ UNA TECLA (SÓLO DURA UN CICLO DE RELOJ)
	);

END LIB_TEC_MATRICIAL_4x4_INTESC_RevA;

ARCHITECTURE Behavioral OF LIB_TEC_MATRICIAL_4x4_INTESC_RevA IS

	CONSTANT DELAY_1MS : INTEGER := (FREQ_CLK/1000) - 1;
	CONSTANT DELAY_10MS : INTEGER := (FREQ_CLK/100) - 1;

	SIGNAL CONTA_1MS : INTEGER RANGE 0 TO DELAY_1MS := 0;
	SIGNAL BANDERA : STD_LOGIC := '0';
	SIGNAL CONTA_10MS : INTEGER RANGE 0 TO DELAY_10MS := 0;
	SIGNAL BANDERA2 : STD_LOGIC := '0';

	SIGNAL REG_B1 : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL REG_B2 : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL REG_B3 : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL REG_B4 : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL REG_B5 : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL REG_B6 : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL REG_B7 : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL REG_B8 : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL REG_B9 : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL REG_BA : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL REG_BB : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL REG_BC : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL REG_BD : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL REG_B0 : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL REG_BAS : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');
	SIGNAL REG_BGA : STD_LOGIC_VECTOR(7 DOWNTO 0) := (OTHERS => '0');

	SIGNAL FILA_REG_S : STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
	SIGNAL FILA : INTEGER RANGE 0 TO 3 := 0;

	SIGNAL IND_S : STD_LOGIC := '0';
	SIGNAL EDO : INTEGER RANGE 0 TO 1 := 0;

BEGIN

	FILAS <= FILA_REG_S;

	--RETARDO 1 MS--
	PROCESS (CLK)
	BEGIN
		IF RISING_EDGE(CLK) THEN
			CONTA_1MS <= CONTA_1MS + 1;
			BANDERA <= '0';
			IF CONTA_1MS = DELAY_1MS THEN
				CONTA_1MS <= 0;
				BANDERA <= '1';
			END IF;
		END IF;
	END PROCESS;
	----------------

	--RETARDO 10 MS--
	PROCESS (CLK)
	BEGIN
		IF RISING_EDGE(CLK) THEN
			CONTA_10MS <= CONTA_10MS + 1;
			BANDERA2 <= '0';
			IF CONTA_10MS = DELAY_10MS THEN
				CONTA_10MS <= 0;
				BANDERA2 <= '1';
			END IF;
		END IF;
	END PROCESS;
	----------------

	--PROCESO QUE ACTIVA CADA FILA CADA 10ms--
	PROCESS (CLK, BANDERA2)
	BEGIN
		IF RISING_EDGE(CLK) AND BANDERA2 = '1' THEN
			FILA <= FILA + 1;
			IF FILA = 3 THEN
				FILA <= 0;
			END IF;
		END IF;
	END PROCESS;

	WITH FILA SELECT
		FILA_REG_S <= "1000" WHEN 0,
		"0100" WHEN 1,
		"0010" WHEN 2,
		"0001" WHEN OTHERS;
	-------------------------------				

	----------PROCESO QUE EVITA EL EFECTO REBOTE DE LAS TECLAS----------------
	--LLENA LOS REGISTROS CON '1' DEPENDIENDO EL BOTÓN QUE SE HAYA PRESIONADO--
	PROCESS (CLK, BANDERA)
	BEGIN
		IF RISING_EDGE(CLK) AND BANDERA = '1' THEN
			IF FILA_REG_S = "1000" THEN --PRIMERA FILA DE BOTONES
				REG_B1 <= REG_B1(6 DOWNTO 0) & COLUMNAS(3);
				REG_B2 <= REG_B2(6 DOWNTO 0) & COLUMNAS(2);
				REG_B3 <= REG_B3(6 DOWNTO 0) & COLUMNAS(1);
				REG_BA <= REG_BA(6 DOWNTO 0) & COLUMNAS(0);
			ELSIF FILA_REG_S = "0100" THEN --SEGUNDA FILA DE BOTONES
				REG_B4 <= REG_B4(6 DOWNTO 0) & COLUMNAS(3);
				REG_B5 <= REG_B5(6 DOWNTO 0) & COLUMNAS(2);
				REG_B6 <= REG_B6(6 DOWNTO 0) & COLUMNAS(1);
				REG_BB <= REG_BB(6 DOWNTO 0) & COLUMNAS(0);
			ELSIF FILA_REG_S = "0010" THEN --TERCERA FILA DE BOTONES
				REG_B7 <= REG_B7(6 DOWNTO 0) & COLUMNAS(3);
				REG_B8 <= REG_B8(6 DOWNTO 0) & COLUMNAS(2);
				REG_B9 <= REG_B9(6 DOWNTO 0) & COLUMNAS(1);
				REG_BC <= REG_BC(6 DOWNTO 0) & COLUMNAS(0);
			ELSIF FILA_REG_S = "0001" THEN --CUARTA FILA DE BOTONES
				REG_BAS <= REG_BAS(6 DOWNTO 0) & COLUMNAS(3);
				REG_B0 <= REG_B0(6 DOWNTO 0) & COLUMNAS(2);
				REG_BGA <= REG_BGA(6 DOWNTO 0) & COLUMNAS(1);
				REG_BD <= REG_BD(6 DOWNTO 0) & COLUMNAS(0);
			END IF;
		END IF;
	END PROCESS;
	----------------------------------------------------------------------------

	--MANDA EL DATO A LA SALIDA--
	PROCESS (CLK)
	BEGIN
		IF RISING_EDGE(CLK) THEN
			IF REG_B0 = "11111111" THEN
				BOTON_PRES <= X"0";
				IND_S <= '1';
			ELSIF REG_B1 = "11111111" THEN
				BOTON_PRES <= X"1";
				IND_S <= '1';
			ELSIF REG_B2 = "11111111" THEN
				BOTON_PRES <= X"2";
				IND_S <= '1';
			ELSIF REG_B3 = "11111111" THEN
				BOTON_PRES <= X"3";
				IND_S <= '1';
			ELSIF REG_B4 = "11111111" THEN
				BOTON_PRES <= X"4";
				IND_S <= '1';
			ELSIF REG_B5 = "11111111" THEN
				BOTON_PRES <= X"5";
				IND_S <= '1';
			ELSIF REG_B6 = "11111111" THEN
				BOTON_PRES <= X"6";
				IND_S <= '1';
			ELSIF REG_B7 = "11111111" THEN
				BOTON_PRES <= X"7";
				IND_S <= '1';
			ELSIF REG_B8 = "11111111" THEN
				BOTON_PRES <= X"8";
				IND_S <= '1';
			ELSIF REG_B9 = "11111111" THEN
				BOTON_PRES <= X"9";
				IND_S <= '1';
			ELSIF REG_BA = "11111111" THEN
				BOTON_PRES <= X"A";
				IND_S <= '1';
			ELSIF REG_BB = "11111111" THEN
				BOTON_PRES <= X"B";
				IND_S <= '1';
			ELSIF REG_BC = "11111111" THEN
				BOTON_PRES <= X"C";
				IND_S <= '1';
			ELSIF REG_BD = "11111111" THEN
				BOTON_PRES <= X"D";
				IND_S <= '1';
			ELSIF REG_BAS = "11111111" THEN
				BOTON_PRES <= X"E";
				IND_S <= '1';
			ELSIF REG_BGA = "11111111" THEN
				BOTON_PRES <= X"F";
				IND_S <= '1';
			ELSE
				IND_S <= '0';
			END IF;
		END IF;
	END PROCESS;
	-----------------------------

	--MÁQUINA DE ESTADOS PARA LA BANDERA--
	PROCESS (CLK)
	BEGIN
		IF RISING_EDGE(CLK) THEN
			IF EDO = 0 THEN
				IF IND_S = '1' THEN
					IND <= '1';
					EDO <= 1;
				ELSE
					EDO <= 0;
					IND <= '0';
				END IF;
			ELSE
				IF IND_S = '1' THEN
					EDO <= 1;
					IND <= '0';
				ELSE
					EDO <= 0;
				END IF;
			END IF;
		END IF;
	END PROCESS;
	--------------------------------------
END Behavioral;